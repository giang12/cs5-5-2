
module xor2_47 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_46 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_15 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_45 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_44 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_43 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_14 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_42 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_41 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_40 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_13 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_39 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_38 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_37 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_12 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_36 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_35 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_34 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_11 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_33 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_32 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_31 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_10 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_30 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_29 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_28 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_9 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_27 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_26 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_25 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_8 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_24 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_23 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_22 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_7 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_21 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_20 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_19 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_6 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_18 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_17 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_16 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_5 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_15 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_14 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_13 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_4 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_12 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_11 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_10 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_3 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_9 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_8 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_7 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_2 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_6 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_5 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_4 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_1 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_3 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_2 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_1 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module and2_0 ( out, in1, in2 );
  input in1, in2;
  output out;


  AND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_0 ( out, in1, in2 );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module fulladder_15 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_47 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_46 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_15 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_45 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_14 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_44 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_43 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_14 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_42 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_13 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_41 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_40 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_13 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_39 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_12 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_38 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_37 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_12 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_36 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_11 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_35 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_34 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_11 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_33 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_10 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_32 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_31 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_10 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_30 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_9 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_29 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_28 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_9 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_27 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_8 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_26 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_25 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_8 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_24 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_7 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_23 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_22 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_7 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_21 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_6 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_20 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_19 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_6 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_18 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_5 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_17 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_16 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_5 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_15 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_4 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_14 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_13 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_4 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_12 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_3 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_11 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_10 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_3 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_9 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_2 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_8 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_7 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_2 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_6 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_1 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_5 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_4 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_1 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_3 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_0 ( S, P, G, InA, InB, Cin );
  input InA, InB, Cin;
  output S, P, G;
  wire   w1;

  xor2_2 mod1 ( .out(w1), .in1(InB), .in2(Cin) );
  xor2_1 mod2 ( .out(S), .in1(InA), .in2(w1) );
  and2_0 mod3 ( .out(G), .in1(InA), .in2(InB) );
  xor2_0 mod4 ( .out(P), .in1(InA), .in2(InB) );
endmodule


module fulladder_16bit ( .S({\S<15> , \S<14> , \S<13> , \S<12> , \S<11> , 
        \S<10> , \S<9> , \S<8> , \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , 
        \S<2> , \S<1> , \S<0> }), .P({\P<15> , \P<14> , \P<13> , \P<12> , 
        \P<11> , \P<10> , \P<9> , \P<8> , \P<7> , \P<6> , \P<5> , \P<4> , 
        \P<3> , \P<2> , \P<1> , \P<0> }), .G({\G<15> , \G<14> , \G<13> , 
        \G<12> , \G<11> , \G<10> , \G<9> , \G<8> , \G<7> , \G<6> , \G<5> , 
        \G<4> , \G<3> , \G<2> , \G<1> , \G<0> }), .A({\A<15> , \A<14> , 
        \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> , \A<7> , \A<6> , 
        \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<15> , \B<14> , 
        \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> , \B<7> , \B<6> , 
        \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> }), .CI({\CI<15> , 
        \CI<14> , \CI<13> , \CI<12> , \CI<11> , \CI<10> , \CI<9> , \CI<8> , 
        \CI<7> , \CI<6> , \CI<5> , \CI<4> , \CI<3> , \CI<2> , \CI<1> , \CI<0> 
        }) );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> ,
         \CI<15> , \CI<14> , \CI<13> , \CI<12> , \CI<11> , \CI<10> , \CI<9> ,
         \CI<8> , \CI<7> , \CI<6> , \CI<5> , \CI<4> , \CI<3> , \CI<2> ,
         \CI<1> , \CI<0> ;
  output \S<15> , \S<14> , \S<13> , \S<12> , \S<11> , \S<10> , \S<9> , \S<8> ,
         \S<7> , \S<6> , \S<5> , \S<4> , \S<3> , \S<2> , \S<1> , \S<0> ,
         \P<15> , \P<14> , \P<13> , \P<12> , \P<11> , \P<10> , \P<9> , \P<8> ,
         \P<7> , \P<6> , \P<5> , \P<4> , \P<3> , \P<2> , \P<1> , \P<0> ,
         \G<15> , \G<14> , \G<13> , \G<12> , \G<11> , \G<10> , \G<9> , \G<8> ,
         \G<7> , \G<6> , \G<5> , \G<4> , \G<3> , \G<2> , \G<1> , \G<0> ;


  fulladder_15 fulladder0 ( .S(\S<0> ), .P(\P<0> ), .G(\G<0> ), .InA(\A<0> ), 
        .InB(\B<0> ), .Cin(\CI<0> ) );
  fulladder_14 fulladder1 ( .S(\S<1> ), .P(\P<1> ), .G(\G<1> ), .InA(\A<1> ), 
        .InB(\B<1> ), .Cin(\CI<1> ) );
  fulladder_13 fulladder2 ( .S(\S<2> ), .P(\P<2> ), .G(\G<2> ), .InA(\A<2> ), 
        .InB(\B<2> ), .Cin(\CI<2> ) );
  fulladder_12 fulladder3 ( .S(\S<3> ), .P(\P<3> ), .G(\G<3> ), .InA(\A<3> ), 
        .InB(\B<3> ), .Cin(\CI<3> ) );
  fulladder_11 fulladder4 ( .S(\S<4> ), .P(\P<4> ), .G(\G<4> ), .InA(\A<4> ), 
        .InB(\B<4> ), .Cin(\CI<4> ) );
  fulladder_10 fulladder5 ( .S(\S<5> ), .P(\P<5> ), .G(\G<5> ), .InA(\A<5> ), 
        .InB(\B<5> ), .Cin(\CI<5> ) );
  fulladder_9 fulladder6 ( .S(\S<6> ), .P(\P<6> ), .G(\G<6> ), .InA(\A<6> ), 
        .InB(\B<6> ), .Cin(\CI<6> ) );
  fulladder_8 fulladder7 ( .S(\S<7> ), .P(\P<7> ), .G(\G<7> ), .InA(\A<7> ), 
        .InB(\B<7> ), .Cin(\CI<7> ) );
  fulladder_7 fulladder8 ( .S(\S<8> ), .P(\P<8> ), .G(\G<8> ), .InA(\A<8> ), 
        .InB(\B<8> ), .Cin(\CI<8> ) );
  fulladder_6 fulladder9 ( .S(\S<9> ), .P(\P<9> ), .G(\G<9> ), .InA(\A<9> ), 
        .InB(\B<9> ), .Cin(\CI<9> ) );
  fulladder_5 fulladder10 ( .S(\S<10> ), .P(\P<10> ), .G(\G<10> ), .InA(
        \A<10> ), .InB(\B<10> ), .Cin(\CI<10> ) );
  fulladder_4 fulladder11 ( .S(\S<11> ), .P(\P<11> ), .G(\G<11> ), .InA(
        \A<11> ), .InB(\B<11> ), .Cin(\CI<11> ) );
  fulladder_3 fulladder12 ( .S(\S<12> ), .P(\P<12> ), .G(\G<12> ), .InA(
        \A<12> ), .InB(\B<12> ), .Cin(\CI<12> ) );
  fulladder_2 fulladder13 ( .S(\S<13> ), .P(\P<13> ), .G(\G<13> ), .InA(
        \A<13> ), .InB(\B<13> ), .Cin(\CI<13> ) );
  fulladder_1 fulladder14 ( .S(\S<14> ), .P(\P<14> ), .G(\G<14> ), .InA(
        \A<14> ), .InB(\B<14> ), .Cin(\CI<14> ) );
  fulladder_0 fulladder15 ( .S(\S<15> ), .P(\P<15> ), .G(\G<15> ), .InA(
        \A<15> ), .InB(\B<15> ), .Cin(\CI<15> ) );
endmodule

