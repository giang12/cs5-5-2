module branch_cond_test(readData1, readData2, IFID_instr, branch, jump, pcSrc);
    input [15:0] readData1, readData2;
    input [1:0] IFID_instr; // IF/ID_instr[12:11]
    input branch, jump;
    output pcSrc;
    
    // your facny code goes here

endmodule
