library verilog;
use verilog.vl_types.all;
entity dff_8bit_tb is
end dff_8bit_tb;
