module cla_4bit (CO, PG, GG, CI, P, G);
    input [3:0] P, G;
    input CI;
    output [3:0] CO;
    output PG, GG;



