module hazard_detect(pcWriteEn, IFIDWriteEn, control_sel, IDEX_Instr, IFID_Instr, IDEX_Mem_En, IDEX_Mem_Wr);

    input [15:0] IDEX_Instr, IFID_Instr;
    input IDEX_Mem_En, IDEX_Mem_Wr;
    output pcWriteEn, IFIDWriteEn, control_sel;

    // your fancy code goes here
    

endmodule
