library verilog;
use verilog.vl_types.all;
entity dff_16bit_tb is
end dff_16bit_tb;
