module forward_unit(ALUSel1, ALUSel2, IDEX_Instr, EXMEM_Instr, MEMWB_Instr, EXMEM_wb, MEMWB_wb); 
    input [15:0] IDEX_Instr, EXMEM_Instr, MEMWB_Instr;
    input EXMEM_wb, MEMWB_wb;
    output ALUSel1, ALUSel2;
    
    // your fancy code goes here
    

    
endmodule

