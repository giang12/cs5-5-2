module regEXMem();
    input 
    output

    // Control Portion
    

    // Data Portion


endmodule

