module regIFID();
    input 
    output

    // Control Portion
    

    // Data Portion


endmodule

