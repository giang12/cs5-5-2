module regMemWB();
    input 
    output

    // Control Portion
    

    // Data Portion


endmodule

