module cla_4bit(P, G, CI, CO);
input [3:0] P, G;
input CI;
output [3:0] CO;
output PG, GG;


