module regIDEX();
    input 
    output

    // Control Portion
    

    // Data Portion


endmodule

