library verilog;
use verilog.vl_types.all;
entity reg_64bit_tb is
end reg_64bit_tb;
