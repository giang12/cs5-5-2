module and3(out, in1, in2, in3);
input in1, in2, in3;
output out;
assign out = in1 & in2 & in3;
endmodule
