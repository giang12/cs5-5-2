module cond_set(cond, instr, zero, Ofl, out);
    input zero, Ofl, out;
    input [1:0] instr;
    output [15:0] cond;


endmodule
